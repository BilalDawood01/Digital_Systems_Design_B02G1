LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY x2sin IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      x        :  IN    STD_LOGIC_VECTOR(8 DOWNTO 0);                           
      sinx       :  OUT   STD_LOGIC_VECTOR(8 DOWNTO 0));  
END x2sin;

ARCHITECTURE behavior OF x2sin IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are duty cycles. They are determined via
-- the following formula: (511/2) * (sin(x)+1). 511 = 2^(9) - 1.
-- The indexes are x values. 

type array_1d is array (0 to 511) of integer;
constant x2s_LUT : array_1d := (


( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 1 ) ,
( 1 ) ,
( 1 ) ,
( 2 ) ,
( 2 ) ,
( 3 ) ,
( 3 ) ,
( 4 ) ,
( 4 ) ,
( 5 ) ,
( 6 ) ,
( 6 ) ,
( 7 ) ,
( 8 ) ,
( 9 ) ,
( 10 ) ,
( 11 ) ,
( 11 ) ,
( 12 ) ,
( 13 ) ,
( 14 ) ,
( 16 ) ,
( 17 ) ,
( 18 ) ,
( 19 ) ,
( 20 ) ,
( 21 ) ,
( 23 ) ,
( 24 ) ,
( 25 ) ,
( 27 ) ,
( 28 ) ,
( 30 ) ,
( 31 ) ,
( 33 ) ,
( 34 ) ,
( 36 ) ,
( 38 ) ,
( 39 ) ,
( 41 ) ,
( 43 ) ,
( 44 ) ,
( 46 ) ,
( 48 ) ,
( 50 ) ,
( 52 ) ,
( 54 ) ,
( 56 ) ,
( 58 ) ,
( 60 ) ,
( 62 ) ,
( 64 ) ,
( 66 ) ,
( 68 ) ,
( 70 ) ,
( 72 ) ,
( 74 ) ,
( 77 ) ,
( 79 ) ,
( 81 ) ,
( 84 ) ,
( 86 ) ,
( 88 ) ,
( 91 ) ,
( 93 ) ,
( 96 ) ,
( 98 ) ,
( 100 ) ,
( 103 ) ,
( 106 ) ,
( 108 ) ,
( 111 ) ,
( 113 ) ,
( 116 ) ,
( 119 ) ,
( 121 ) ,
( 124 ) ,
( 127 ) ,
( 129 ) ,
( 132 ) ,
( 135 ) ,
( 138 ) ,
( 140 ) ,
( 143 ) ,
( 146 ) ,
( 149 ) ,
( 152 ) ,
( 155 ) ,
( 157 ) ,
( 160 ) ,
( 163 ) ,
( 166 ) ,
( 169 ) ,
( 172 ) ,
( 175 ) ,
( 178 ) ,
( 181 ) ,
( 184 ) ,
( 187 ) ,
( 190 ) ,
( 193 ) ,
( 196 ) ,
( 199 ) ,
( 202 ) ,
( 206 ) ,
( 209 ) ,
( 212 ) ,
( 215 ) ,
( 218 ) ,
( 221 ) ,
( 224 ) ,
( 227 ) ,
( 230 ) ,
( 233 ) ,
( 237 ) ,
( 240 ) ,
( 243 ) ,
( 246 ) ,
( 249 ) ,
( 252 ) ,
( 256 ) ,
( 259 ) ,
( 262 ) ,
( 265 ) ,
( 268 ) ,
( 271 ) ,
( 274 ) ,
( 277 ) ,
( 281 ) ,
( 284 ) ,
( 287 ) ,
( 290 ) ,
( 293 ) ,
( 296 ) ,
( 299 ) ,
( 302 ) ,
( 305 ) ,
( 309 ) ,
( 312 ) ,
( 315 ) ,
( 318 ) ,
( 321 ) ,
( 324 ) ,
( 327 ) ,
( 330 ) ,
( 333 ) ,
( 336 ) ,
( 339 ) ,
( 342 ) ,
( 345 ) ,
( 348 ) ,
( 351 ) ,
( 353 ) ,
( 356 ) ,
( 359 ) ,
( 362 ) ,
( 365 ) ,
( 368 ) ,
( 371 ) ,
( 373 ) ,
( 376 ) ,
( 379 ) ,
( 382 ) ,
( 384 ) ,
( 387 ) ,
( 390 ) ,
( 392 ) ,
( 395 ) ,
( 398 ) ,
( 400 ) ,
( 403 ) ,
( 405 ) ,
( 408 ) ,
( 411 ) ,
( 413 ) ,
( 415 ) ,
( 418 ) ,
( 420 ) ,
( 423 ) ,
( 425 ) ,
( 427 ) ,
( 430 ) ,
( 432 ) ,
( 434 ) ,
( 437 ) ,
( 439 ) ,
( 441 ) ,
( 443 ) ,
( 445 ) ,
( 447 ) ,
( 449 ) ,
( 451 ) ,
( 453 ) ,
( 455 ) ,
( 457 ) ,
( 459 ) ,
( 461 ) ,
( 463 ) ,
( 465 ) ,
( 467 ) ,
( 468 ) ,
( 470 ) ,
( 472 ) ,
( 473 ) ,
( 475 ) ,
( 477 ) ,
( 478 ) ,
( 480 ) ,
( 481 ) ,
( 483 ) ,
( 484 ) ,
( 486 ) ,
( 487 ) ,
( 488 ) ,
( 490 ) ,
( 491 ) ,
( 492 ) ,
( 493 ) ,
( 494 ) ,
( 495 ) ,
( 497 ) ,
( 498 ) ,
( 499 ) ,
( 500 ) ,
( 500 ) ,
( 501 ) ,
( 502 ) ,
( 503 ) ,
( 504 ) ,
( 505 ) ,
( 505 ) ,
( 506 ) ,
( 507 ) ,
( 507 ) ,
( 508 ) ,
( 508 ) ,
( 509 ) ,
( 509 ) ,
( 510 ) ,
( 510 ) ,
( 510 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 510 ) ,
( 510 ) ,
( 510 ) ,
( 509 ) ,
( 509 ) ,
( 508 ) ,
( 508 ) ,
( 507 ) ,
( 507 ) ,
( 506 ) ,
( 505 ) ,
( 505 ) ,
( 504 ) ,
( 503 ) ,
( 502 ) ,
( 501 ) ,
( 500 ) ,
( 500 ) ,
( 499 ) ,
( 498 ) ,
( 497 ) ,
( 495 ) ,
( 494 ) ,
( 493 ) ,
( 492 ) ,
( 491 ) ,
( 490 ) ,
( 488 ) ,
( 487 ) ,
( 486 ) ,
( 484 ) ,
( 483 ) ,
( 481 ) ,
( 480 ) ,
( 478 ) ,
( 477 ) ,
( 475 ) ,
( 473 ) ,
( 472 ) ,
( 470 ) ,
( 468 ) ,
( 467 ) ,
( 465 ) ,
( 463 ) ,
( 461 ) ,
( 459 ) ,
( 457 ) ,
( 455 ) ,
( 453 ) ,
( 451 ) ,
( 449 ) ,
( 447 ) ,
( 445 ) ,
( 443 ) ,
( 441 ) ,
( 439 ) ,
( 437 ) ,
( 434 ) ,
( 432 ) ,
( 430 ) ,
( 427 ) ,
( 425 ) ,
( 423 ) ,
( 420 ) ,
( 418 ) ,
( 415 ) ,
( 413 ) ,
( 411 ) ,
( 408 ) ,
( 405 ) ,
( 403 ) ,
( 400 ) ,
( 398 ) ,
( 395 ) ,
( 392 ) ,
( 390 ) ,
( 387 ) ,
( 384 ) ,
( 382 ) ,
( 379 ) ,
( 376 ) ,
( 373 ) ,
( 371 ) ,
( 368 ) ,
( 365 ) ,
( 362 ) ,
( 359 ) ,
( 356 ) ,
( 353 ) ,
( 351 ) ,
( 348 ) ,
( 345 ) ,
( 342 ) ,
( 339 ) ,
( 336 ) ,
( 333 ) ,
( 330 ) ,
( 327 ) ,
( 324 ) ,
( 321 ) ,
( 318 ) ,
( 315 ) ,
( 312 ) ,
( 309 ) ,
( 305 ) ,
( 302 ) ,
( 299 ) ,
( 296 ) ,
( 293 ) ,
( 290 ) ,
( 287 ) ,
( 284 ) ,
( 281 ) ,
( 277 ) ,
( 274 ) ,
( 271 ) ,
( 268 ) ,
( 265 ) ,
( 262 ) ,
( 259 ) ,
( 256 ) ,
( 252 ) ,
( 249 ) ,
( 246 ) ,
( 243 ) ,
( 240 ) ,
( 237 ) ,
( 234 ) ,
( 230 ) ,
( 227 ) ,
( 224 ) ,
( 221 ) ,
( 218 ) ,
( 215 ) ,
( 212 ) ,
( 209 ) ,
( 206 ) ,
( 203 ) ,
( 199 ) ,
( 196 ) ,
( 193 ) ,
( 190 ) ,
( 187 ) ,
( 184 ) ,
( 181 ) ,
( 178 ) ,
( 175 ) ,
( 172 ) ,
( 169 ) ,
( 166 ) ,
( 163 ) ,
( 160 ) ,
( 158 ) ,
( 155 ) ,
( 152 ) ,
( 149 ) ,
( 146 ) ,
( 143 ) ,
( 140 ) ,
( 138 ) ,
( 135 ) ,
( 132 ) ,
( 129 ) ,
( 127 ) ,
( 124 ) ,
( 121 ) ,
( 119 ) ,
( 116 ) ,
( 113 ) ,
( 111 ) ,
( 108 ) ,
( 106 ) ,
( 103 ) ,
( 101 ) ,
( 98 ) ,
( 96 ) ,
( 93 ) ,
( 91 ) ,
( 88 ) ,
( 86 ) ,
( 84 ) ,
( 81 ) ,
( 79 ) ,
( 77 ) ,
( 75 ) ,
( 72 ) ,
( 70 ) ,
( 68 ) ,
( 66 ) ,
( 64 ) ,
( 62 ) ,
( 60 ) ,
( 58 ) ,
( 56 ) ,
( 54 ) ,
( 52 ) ,
( 50 ) ,
( 48 ) ,
( 46 ) ,
( 44 ) ,
( 43 ) ,
( 41 ) ,
( 39 ) ,
( 38 ) ,
( 36 ) ,
( 34 ) ,
( 33 ) ,
( 31 ) ,
( 30 ) ,
( 28 ) ,
( 27 ) ,
( 25 ) ,
( 24 ) ,
( 23 ) ,
( 21 ) ,
( 20 ) ,
( 19 ) ,
( 18 ) ,
( 17 ) ,
( 16 ) ,
( 14 ) ,
( 13 ) ,
( 12 ) ,
( 11 ) ,
( 11 ) ,
( 10 ) ,
( 9 ) ,
( 8 ) ,
( 7 ) ,
( 6 ) ,
( 6 ) ,
( 5 ) ,
( 4 ) ,
( 4 ) ,
( 3 ) ,
( 3 ) ,
( 2 ) ,
( 2 ) ,
( 1 ) ,
( 1 ) ,
( 1 ) 

);


begin
    	
   sinx <= std_logic_vector(to_unsigned(x2s_LUT(to_integer(unsigned(x))),sinx'length));

end behavior;
