LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY x2square IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      x        :  IN    STD_LOGIC_VECTOR(11 DOWNTO 0);                           
      sinx       :  OUT   STD_LOGIC_VECTOR(8 DOWNTO 0));  
END x2square;

ARCHITECTURE behavior OF x2square IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are duty cycles. They are determined via
-- the following formula: (511/2) * (sin(x)+1). 511 = 2^(9) - 1.
-- The indexes are x values. 

type array_1d is array (0 to 4095) of integer;
constant x2s_LUT : array_1d := (

( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 0 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) ,
( 511 ) 



);


begin
    	
   sinx <= std_logic_vector(to_unsigned(x2s_LUT(to_integer(unsigned(x))),sinx'length));

end behavior;
